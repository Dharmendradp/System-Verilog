class base_pkt;
randc bit [1:0]Din;
bit rst;
bit [1:0]Q;
endclass :base_pkt


