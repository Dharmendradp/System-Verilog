package env_package;

`include "base_pkt.sv";
`include "driver.sv";
`include "generator.sv";
`include "monitor.sv";
`include "scoreboard.sv";

endpackage :env_package
